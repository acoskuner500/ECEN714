/home/grads/a/acoskuner500/cadence/synthesis/cru_con/iit018_stdcells.lef